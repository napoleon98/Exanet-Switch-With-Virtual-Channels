`timescale 1ns / 1ps
import exanet_crosb_pkg::*;
import exanet_pkg::*;



module exa_crosb_e2s_with_VCs_tb(

);
  
  localparam prio_num = 2;
  localparam vc_num = 3;
  localparam output_num = 8;
  
  
  reg                     clk		    = 0;
  always #5 clk = ~clk;
  reg                     resetn	    = 0;


  
  exanet s_exanet_tx();   
  AXIS m_axis();  
  reg  traffic_work;
  reg [2:0] rand_2 = 0;
  reg [2:0] rand_3 = 0;

  reg [5:0] rand_6 = 0;
  logic [4:0] header_vc;
  cntrl_info_t                  cntrl_info;
  

  //each traffic generator creates a file, and writes in it, the various details 
  //of each packet generated by it. (the packet is randomly generated). it then
  //"tags" the address of this packet on the "CRC" part of the header which is not
  //used by the switch    
  exa_crosb_traffic_gen #(
          .tag(0),
          .vc_num(vc_num)
     )traffic_gen_0 (
          .clk(clk),
          .resetn(resetn),
          .i_src_coord(0),
          .dif_size_enable(0),
          .dif_type_enable(0),
          .fixed_dest_enable(1),//it was 1
          .fixed_header_vc_enable(0),
          .fixed_dest(0),//10
          .i_work(traffic_work),
          .exa(s_exanet_tx),
          .valid_drop_rate(0),
          .fixed_header_vc(0)
        ); 
        
         
   
   
   
 
  
    
  logic [prio_num*vc_num-1 : 0] has_packet; 
  
  logic [prio_num*vc_num-1 : 0] fifo_full;
  logic [output_num-1 : 0] out_fifo_credits [vc_num-1 : 0];
  logic [vc_num-1 :0] high_prio_requests;
  logic [vc_num-1 :0] low_prio_requests;
  logic [$clog2(output_num)-1 :0]  dests[prio_num*vc_num-1 : 0] ;
  //outputs
  logic [prio_num*vc_num- 1: 0] selected_vc_from_input_arbiter;  
  logic cts_from_input_arbiter;
   
  exa_crosb_e2s_with_VCs # (
         .fifo_enable          (1),
         .prio_num             (prio_num),
         .vc_num               (vc_num),
         .net_route_reg_enable (0),
         .in_fifo_depth        (64),
         .TDEST_WIDTH          (),
         .output_num           (output_num),
         .max_ports            (8),
         .PORTx_LOW_ADDR   ({42'h38000000000,42'h38000000010,42'h38000000020,42'h38000000030,42'h38000000040,42'h38000000050,42'h38000000060,42'h38000000070} ),//{42'h38000000000}
         .PORTx_HIGH_ADDR  ({42'h38000000010,42'h38000000020,42'h38000000030,42'h38000000040,42'h38000000050,42'h38000000060,42'h38000000070,42'h38000000080} )//{42'h380000fffff}
     ) e2s_dut   (
            // AXI STREAM IF
         .M_ACLK(clk),
         .M_ARESETN(resetn),
         .i_src_coord(0),
         .M_AXIS(m_axis),    
         .exanet_rx(s_exanet_tx),
         .i_cntrl_info('b0),
         .i_cts_from_input_arbiter(cts_from_input_arbiter),//added
         .i_selected_vc_from_input_arbiter(selected_vc_from_input_arbiter),//added
         .o_dec_error(),
         .o_pkt_counter(),
         .o_has_packet(has_packet),
         .o_fifo_full(fifo_full),
         .o_dests(dests) // added
       ); 
  
  task cts (input [prio_num*vc_num-1:0] selected_vc ); begin
    //#210
    /*
    while(!has_packet[selected_vc]) @(posedge clk);
    @(negedge clk);
     */ 
    selected_vc_from_input_arbiter = selected_vc; 
    cts_from_input_arbiter         = 1;
      
      
    while(!m_axis.TLAST) @(posedge clk); 
    @(negedge clk);
      
    cts_from_input_arbiter           = 0;
  end
  endtask
  
       
  initial begin
    m_axis.TREADY                  = 0;
    traffic_work                   = 0; 
    selected_vc_from_input_arbiter = 0;
    cts_from_input_arbiter         = 0;
    header_vc                      = 0;
    
    #100
    resetn                         = 1;
   
    #100
    traffic_work                   = 1;
    /*
    while(header_vc<6) begin
      while(!fifo_full[header_vc]) @(posedge clk);
      @(negedge clk);
      header_vc                      = header_vc + 1;
      */
     
     while(!fifo_full[0]) begin
       
       @(posedge clk);
     end
       
    
   
  end
  
  
  
  initial begin
   
   rand_6 = $urandom() % 20 + 40 ;
   repeat(rand_6) @(posedge clk);
   
   forever begin
     if(has_packet != 0) begin 
     
       rand_2 = $urandom() % 6;
       while(!has_packet[rand_2]) begin
         rand_2 = $urandom() % 6;
       end
     
       cts(rand_2);
     
       repeat(rand_6) @(posedge clk);
     end   
   end
   
   
    
    
  end


    
endmodule
