`define log2(x) \
 (x >= 1 && x <= 2) ? 1 : \
 (x >= 3 && x <= 4) ? 2 : \
 (x >= 5 && x <= 8) ? 3 : \
 (x >= 9 && x <= 16) ? 4 : \
 (x >= 17 && x <= 32) ? 5 : \
 (x >= 33 && x <= 64) ? 6 : \
 (x >= 65 && x <= 128) ? 7 : \
 (x >= 129 && x <= 256) ? 8 : \
 (x >= 257 && x <= 512) ? 9 : \
 (x >= 513 && x <= 1024) ? 10 : \
 (x >= 1025 && x <= 2048) ? 11 : \
 (x >= 2049 && x <= 4096) ? 12 : \
 (x >= 4097 && x <= 8192) ? 13 : \
 (x >= 8193 && x <= 16384) ? 14 : \
 (x >= 16385 && x <= 32768) ? 15 : \
 (x >= 32769 && x <= 65536) ? 16 : \
 (x >= 65537 && x <= 131072) ? 17 : \
 -1